0.8377202
0
0
0
0
0
0
0
0
0
0